11f7a98aa2eb573689b6ec06123a2df9f2a0b7b2